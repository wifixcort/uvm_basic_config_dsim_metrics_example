`include "uvm_macros.svh"
import uvm_pkg::*;

interface arb_intf(input logic clk);
  
 

endinterface
