`include "uvm_macros.svh"
import uvm_pkg::*;


// `include "../testbench/top_hvl.sv"
`include "../testbench/interface.sv"
`include "../testbench/driver.sv"
`include "../testbench/env.sv"
`include "../testbench/test_basic.sv"
