`include "../rtl/arbiter.v"
`include "../rtl/top_hdl.sv"
